module sine(degrees, d1, d2, d3, d4);  // Просто обрабатываем 360 кейсов
	input [13:0] degrees;
	output reg [7:0] d1;
	output reg [7:0] d2;
	output reg [7:0] d3;
	output reg [7:0] d4;
	always @(degrees) begin
	case (degrees)
	0: begin
    		d1 = 8'b00000001;
    		d2 = 8'b10000001;
    		d3 = 8'b10000001;
    		d4 = 8'b10000001;
    		end
	1: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b11001111;
	    d4 = 8'b10001111;
	    end
	2: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10000110;
	    d4 = 8'b10100100;
	    end
	3: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10100100;
	    d4 = 8'b10010010;
	    end
	4: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	5: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10000000;
	    d4 = 8'b10001111;
	    end
	6: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10100100;
	    end
	7: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10010010;
	    d4 = 8'b10010010;
	    end
	8: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	9: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	10: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	11: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	12: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10000001;
	    d4 = 8'b10000000;
	    end
	13: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10010010;
	    d4 = 8'b10100100;
	    end
	14: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	15: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	16: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10001111;
	    d4 = 8'b10100000;
	    end
	17: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10000100;
	    d4 = 8'b10010010;
	    end
	18: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	19: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10010010;
	    d4 = 8'b10100000;
	    end
	20: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	21: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10100100;
	    d4 = 8'b10000000;
	    end
	22: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	23: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	24: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	25: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10010010;
	    d4 = 8'b10000110;
	    end
	26: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000000;
	    end
	27: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001100;
	    end
	28: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	29: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	30: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10000001;
	    d4 = 8'b10000001;
	    end
	31: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b11001111;
	    d4 = 8'b10100100;
	    end
	32: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000001;
	    end
	33: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100100;
	    end
	34: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	35: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	36: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	37: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10000001;
	    d4 = 8'b10010010;
	    end
	38: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b11001111;
	    d4 = 8'b10100000;
	    end
	39: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	40: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	41: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	42: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	43: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	44: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	45: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	46: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	47: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000110;
	    d4 = 8'b11001111;
	    end
	48: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	49: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100100;
	    end
	50: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	51: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10001111;
	    d4 = 8'b10001111;
	    end
	52: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	53: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	54: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	55: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	56: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	57: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	58: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000000;
	    end
	59: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10100100;
	    d4 = 8'b10001111;
	    end
	60: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	61: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	62: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000000;
	    d4 = 8'b10000110;
	    end
	63: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	64: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	65: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000001;
	    d4 = 8'b10100000;
	    end
	66: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b11001111;
	    d4 = 8'b11001100;
	    end
	67: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b11001111;
	    end
	68: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b10001111;
	    end
	69: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000110;
	    d4 = 8'b11001100;
	    end
	70: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10000001;
	    end
	71: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100000;
	    end
	72: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001111;
	    end
	73: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	74: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b11001111;
	    end
	75: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	76: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	77: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	78: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000000;
	    end
	79: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	80: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	81: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	82: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000001;
	    end
	83: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000110;
	    end
	84: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	85: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100000;
	    end
	86: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000000;
	    end
	87: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	88: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	89: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	90: begin
	    d1 = 8'b01001111;
	    d2 = 8'b10000001;
	    d3 = 8'b10000001;
	    d4 = 8'b10000001;
	    end
	91: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	92: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	93: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	94: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000000;
	    end
	95: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100000;
	    end
	96: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	97: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000110;
	    end
	98: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000001;
	    end
	99: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	100: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	101: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	102: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000000;
	    end
	103: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	104: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	105: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	106: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b11001111;
	    end
	107: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	108: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001111;
	    end
	109: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100000;
	    end
	110: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10000001;
	    end
	111: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000110;
	    d4 = 8'b11001100;
	    end
	112: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b10001111;
	    end
	113: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b11001111;
	    end
	114: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b11001111;
	    d4 = 8'b11001100;
	    end
	115: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000100;
	    d3 = 8'b10000001;
	    d4 = 8'b10100000;
	    end
	116: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	117: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	118: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000000;
	    d4 = 8'b10000110;
	    end
	119: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	120: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	121: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10100100;
	    d4 = 8'b10001111;
	    end
	122: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000000;
	    end
	123: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	124: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	125: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	126: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000000;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	127: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	128: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	129: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10001111;
	    d4 = 8'b10001111;
	    end
	130: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	131: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100100;
	    end
	132: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	133: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000110;
	    d4 = 8'b11001111;
	    end
	134: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	135: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	136: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	137: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	138: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	139: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	140: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	141: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	142: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b11001111;
	    d4 = 8'b10100000;
	    end
	143: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100000;
	    d3 = 8'b10000001;
	    d4 = 8'b10010010;
	    end
	144: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	145: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	146: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	147: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100100;
	    end
	148: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000001;
	    end
	149: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b11001111;
	    d4 = 8'b10100100;
	    end
	150: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10100100;
	    d3 = 8'b10000001;
	    d4 = 8'b10000001;
	    end
	151: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	152: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	153: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001100;
	    end
	154: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000000;
	    end
	155: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10010010;
	    d4 = 8'b10000110;
	    end
	156: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001100;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	157: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	158: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	159: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10100100;
	    d4 = 8'b10000000;
	    end
	160: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	161: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10010010;
	    d4 = 8'b10100000;
	    end
	162: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000110;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	163: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10000100;
	    d4 = 8'b10010010;
	    end
	164: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10001111;
	    d4 = 8'b10100000;
	    end
	165: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	166: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	167: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10010010;
	    d4 = 8'b10100100;
	    end
	168: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10010010;
	    d3 = 8'b10000001;
	    d4 = 8'b10000000;
	    end
	169: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	170: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	171: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	172: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	173: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10010010;
	    d4 = 8'b10010010;
	    end
	174: begin
	    d1 = 8'b00000001;
	    d2 = 8'b11001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10100100;
	    end
	175: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10000000;
	    d4 = 8'b10001111;
	    end
	176: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	177: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10100100;
	    d4 = 8'b10010010;
	    end
	178: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10000110;
	    d4 = 8'b10100100;
	    end
	179: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b11001111;
	    d4 = 8'b10001111;
	    end
	180: begin
	    d1 = 8'b00000001;
	    d2 = 8'b10000001;
	    d3 = 8'b10000001;
	    d4 = 8'b10000001;
	    end
	181: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b11001111;
	    d4 = 8'b10001111;
	    end
	182: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10000110;
	    d4 = 8'b10100100;
	    end
	183: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10100100;
	    d4 = 8'b10010010;
	    end
	184: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	185: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10000000;
	    d4 = 8'b10001111;
	    end
	186: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10100100;
	    end
	187: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10010010;
	    d4 = 8'b10010010;
	    end
	188: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	189: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	190: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	191: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	192: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10000001;
	    d4 = 8'b10000000;
	    end
	193: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10010010;
	    d4 = 8'b10100100;
	    end
	194: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	195: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	196: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10001111;
	    d4 = 8'b10100000;
	    end
	197: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10000100;
	    d4 = 8'b10010010;
	    end
	198: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	199: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10010010;
	    d4 = 8'b10100000;
	    end
	200: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	201: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10100100;
	    d4 = 8'b10000000;
	    end
	202: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	203: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	204: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	205: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10010010;
	    d4 = 8'b10000110;
	    end
	206: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000000;
	    end
	207: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001100;
	    end
	208: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	209: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	210: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10000001;
	    d4 = 8'b10000001;
	    end
	211: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b11001111;
	    d4 = 8'b10100100;
	    end
	212: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000001;
	    end
	213: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100100;
	    end
	214: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	215: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	216: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	217: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10000001;
	    d4 = 8'b10010010;
	    end
	218: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b11001111;
	    d4 = 8'b10100000;
	    end
	219: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	220: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	221: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	222: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	223: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	224: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	225: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	226: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	227: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000110;
	    d4 = 8'b11001111;
	    end
	228: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	229: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100100;
	    end
	230: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	231: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10001111;
	    d4 = 8'b10001111;
	    end
	232: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	233: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	234: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	235: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	236: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	237: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	238: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000000;
	    end
	239: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10100100;
	    d4 = 8'b10001111;
	    end
	240: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	241: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	242: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000000;
	    d4 = 8'b10000110;
	    end
	243: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	244: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	245: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000001;
	    d4 = 8'b10100000;
	    end
	246: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b11001111;
	    d4 = 8'b11001100;
	    end
	247: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b11001111;
	    end
	248: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b10001111;
	    end
	249: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000110;
	    d4 = 8'b11001100;
	    end
	250: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10000001;
	    end
	251: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100000;
	    end
	252: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001111;
	    end
	253: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	254: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b11001111;
	    end
	255: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	256: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	257: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	258: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000000;
	    end
	259: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	260: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	261: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	262: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000001;
	    end
	263: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000110;
	    end
	264: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	265: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100000;
	    end
	266: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000000;
	    end
	267: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	268: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	269: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	270: begin
	    d1 = 8'b01001110;
	    d2 = 8'b10000001;
	    d3 = 8'b10000001;
	    d4 = 8'b10000001;
	    end
	271: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	272: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	273: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	274: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000000;
	    end
	275: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100000;
	    end
	276: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	277: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000110;
	    end
	278: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000100;
	    d4 = 8'b10000001;
	    end
	279: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	280: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	281: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	282: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000000;
	    end
	283: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	284: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	285: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	286: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100000;
	    d4 = 8'b11001111;
	    end
	287: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	288: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001111;
	    end
	289: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100000;
	    end
	290: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b11001100;
	    d4 = 8'b10000001;
	    end
	291: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000110;
	    d4 = 8'b11001100;
	    end
	292: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b10001111;
	    end
	293: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10010010;
	    d4 = 8'b11001111;
	    end
	294: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b11001111;
	    d4 = 8'b11001100;
	    end
	295: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000100;
	    d3 = 8'b10000001;
	    d4 = 8'b10100000;
	    end
	296: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	297: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	298: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000000;
	    d4 = 8'b10000110;
	    end
	299: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	300: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	301: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10100100;
	    d4 = 8'b10001111;
	    end
	302: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000000;
	    end
	303: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	304: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	305: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	306: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000000;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	307: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000100;
	    d4 = 8'b10000100;
	    end
	308: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	309: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10001111;
	    d4 = 8'b10001111;
	    end
	310: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10100000;
	    d4 = 8'b10100000;
	    end
	311: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100100;
	    end
	312: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	313: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000110;
	    d4 = 8'b11001111;
	    end
	314: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b11001111;
	    d4 = 8'b10000100;
	    end
	315: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	316: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10000100;
	    d4 = 8'b10100100;
	    end
	317: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10000000;
	    d4 = 8'b10010010;
	    end
	318: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	319: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	320: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b11001100;
	    d4 = 8'b10000110;
	    end
	321: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10010010;
	    d4 = 8'b10000100;
	    end
	322: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b11001111;
	    d4 = 8'b10100000;
	    end
	323: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100000;
	    d3 = 8'b10000001;
	    d4 = 8'b10010010;
	    end
	324: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10000000;
	    d4 = 8'b10000000;
	    end
	325: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	326: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	327: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b11001100;
	    d4 = 8'b10100100;
	    end
	328: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000001;
	    end
	329: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b11001111;
	    d4 = 8'b10100100;
	    end
	330: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10100100;
	    d3 = 8'b10000001;
	    d4 = 8'b10000001;
	    end
	331: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10000000;
	    d4 = 8'b10100100;
	    end
	332: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10100000;
	    d4 = 8'b10000100;
	    end
	333: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10100100;
	    d4 = 8'b11001100;
	    end
	334: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10000110;
	    d4 = 8'b10000000;
	    end
	335: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10010010;
	    d4 = 8'b10000110;
	    end
	336: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001100;
	    d3 = 8'b10000001;
	    d4 = 8'b10001111;
	    end
	337: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	338: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10001111;
	    d4 = 8'b10100100;
	    end
	339: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10100100;
	    d4 = 8'b10000000;
	    end
	340: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	341: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10010010;
	    d4 = 8'b10100000;
	    end
	342: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000110;
	    d3 = 8'b10000001;
	    d4 = 8'b10000100;
	    end
	343: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10000100;
	    d4 = 8'b10010010;
	    end
	344: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10001111;
	    d4 = 8'b10100000;
	    end
	345: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10100100;
	    d4 = 8'b10000100;
	    end
	346: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b11001100;
	    d4 = 8'b10010010;
	    end
	347: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10010010;
	    d4 = 8'b10100100;
	    end
	348: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10010010;
	    d3 = 8'b10000001;
	    d4 = 8'b10000000;
	    end
	349: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10000100;
	    d4 = 8'b11001111;
	    end
	350: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10001111;
	    d4 = 8'b11001100;
	    end
	351: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10100100;
	    d4 = 8'b10100000;
	    end
	352: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10000110;
	    d4 = 8'b10000100;
	    end
	353: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10010010;
	    d4 = 8'b10010010;
	    end
	354: begin
	    d1 = 8'b01111110;
	    d2 = 8'b11001111;
	    d3 = 8'b10000001;
	    d4 = 8'b10100100;
	    end
	355: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10000000;
	    d4 = 8'b10001111;
	    end
	356: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10001111;
	    d4 = 8'b10000001;
	    end
	357: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10100100;
	    d4 = 8'b10010010;
	    end
	358: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b10000110;
	    d4 = 8'b10100100;
	    end
	359: begin
	    d1 = 8'b01111110;
	    d2 = 8'b10000001;
	    d3 = 8'b11001111;
	    d4 = 8'b10001111;
   	    end
	default: begin
		 d1 = 8'b01111110;
	    d2 = 8'b01111110;
	    d3 = 8'b01111110;
	    d4 = 8'b01111110;
			 end
	endcase 
	end
	
endmodule
